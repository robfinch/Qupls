// ============================================================================
//        __
//   \\__/ o\    (C) 2021-2025  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================

import QuplsPkg::*;

module Qupls_decode_load(instr, load, cload, cload_tags);
input instruction_t instr;
output load;
output cload;
output cload_tags;

function fnIsLoad;
input instruction_t op;
begin
	case(op.any.opcode)
	OP_JSRI,
	OP_LDx,OP_FLDx,OP_DFLDx,OP_PLDx,OP_LDxU:
		fnIsLoad = 1'b1;
	default:
		fnIsLoad = 1'b0;
	endcase
end
endfunction

function fnIsCLoad;
input instruction_t op;
begin
	case(op.any.opcode)
	OP_LDCAPx:	fnIsCLoad = 1'b1;
	default:
		fnIsCLoad = 1'b0;
	endcase
end
endfunction

function fnIsCLoadTags;
input instruction_t op;
begin
	case(op.any.opcode)
	OP_CAP:
		case(op.cap.func)
		FN_CLOADTAGS:	fnIsCLoadTags = 1'b1;
		default:	fnIsCLoadTags = 1'b0;
		endcase
	default:
		fnIsCLoadTags = 1'b0;
	endcase
end
endfunction

assign load = fnIsLoad(instr);
assign cload = fnIsCLoad(instr);
assign cload_tags = fnIsCLoad(instr);

endmodule
