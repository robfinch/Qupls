`timescale 1ns / 1ps
// ============================================================================
//        __
//   \\__/ o\    (C) 2026  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================
//

module ht_bounce_counter(rst, clk, max_bounce, xlat, found, vadr, count, cd_vadr);
input rst;
input clk;
input [7:0] max_bounce;
input xlat;
input found;
input [31:0] vadr;
output reg [7:0] count;
output reg cd_vadr;

// Bounce counter

reg [7:0] count1;
reg [31:0] vadr1;
always_ff @(posedge clk)
	vadr1 <= vadr;
always_comb
	if (vadr1 != vadr) begin
		count = 8'd0;
		cd_vadr = TRUE;
	end
	else begin
		count = count1;
		cd_vadr = FALSE;
	end

always_ff @(posedge clk)
if (rst)
	count1 <= 8'd0;
else begin
	if (xlat) begin
		if (!found) begin	// not found
			count1 <= count1 + 8'd1;
			if (count1==max_bounce)
				count1 <= 8'd0;
		end
//		else
//			count1 <= 8'd0;
	end
	if (vadr1 != vadr)
		count1 <= 8'd0;
end

endmodule
