// ============================================================================
//        __
//   \\__/ o\    (C) 2025-2026  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//                        
//	2650 LUTs / 2000 FFs / 7.5 BRAMs
// ============================================================================

import const_pkg::*;
import Qupls4_pkg::*;

module Qupls4_checkpoint_manager(rst, clk, clk5x, ph4, fcu_id,
	mux_hdr_cndx, dec_hdr_cndx, ren_hdr_cndx, pgh,
	setcp, setcp_grp, cndx, freecp, freecp_grp, alloc_chkpt, restore, miss_cp);
parameter MWIDTH = 4;
input rst;
input clk;
input clk5x;
input [4:0] ph4;
input rob_ndx_t fcu_id;
input cpu_types_pkg::checkpt_ndx_t mux_hdr_cndx;
input cpu_types_pkg::checkpt_ndx_t dec_hdr_cndx;
input cpu_types_pkg::checkpt_ndx_t ren_hdr_cndx;
input Qupls4_pkg::pipeline_group_hdr_t [Qupls4_pkg::ROB_ENTRIES/4-1:0] pgh;
output reg setcp;
output reg [5:0] setcp_grp;
output wire freecp;
output wire [5:0] freecp_grp;
output reg alloc_chkpt;

// Checkpoint index. Allocates with a new conditional branch. Future
// instructions will read from the checkpoint files at cndx.
// This is the index used to read the checkpoint RAMs.
// Want the checkpoint to take effect for the next group of instructions.
output cpu_types_pkg::checkpt_ndx_t cndx;
input restore;
input cpu_types_pkg::checkpt_ndx_t miss_cp;

reg ialloc_chkpt;
wire free_chkpt;
assign freecp = free_chkpt;
reg free_chkpt2;
reg [Qupls4_pkg::NCHECK-1:0] chkpts_to_free;
checkpt_ndx_t fchkpt2;
checkpt_ndx_t [3:0] avail_chkpt;
reg [1:0] backout_st2;
reg [5:0] grpcnt;

integer n1;
wire chkpt_stall;
reg [5:0] gndx;
reg [5:0] gndx2;

reg [2:0] wcnt;
always_ff @(posedge clk5x)
if (rst)
	wcnt <= 3'd0;
else begin
	if (ph4[1])
		wcnt <= 3'd0;
	else if (wcnt < 3'd4)
		wcnt <= wcnt + 2'd1;
end

typedef enum logic [1:0] 
{
	CHKPT_IDLE = 2'd0,
	CHKPT_ALLOC1 = 2'd1,
	CHKPT_ALLOC2 = 2'd2,
	CHKPT_SET = 2'd3
} state_t;
state_t state;

// Free all the branch checkpoints no longer in use.
// If it is not used anywhere in the pipeline free it.
always_comb
begin
	chkpts_to_free = {Qupls4_pkg::NCHECK{1'b1}};	// Assume all freeable
	gndx = 6'd0;
	for (gndx = 0; gndx < Qupls4_pkg::ROB_ENTRIES/MWIDTH; gndx = gndx + 1)
		chkpts_to_free[pgh[gndx].cndx] = 1'b0;	// can't free, its being used.
	chkpts_to_free[mux_hdr_cndx] = 1'b0;
	chkpts_to_free[dec_hdr_cndx] = 1'b0;
	chkpts_to_free[ren_hdr_cndx] = 1'b0;
end

// Set checkpoint index
// Backup the checkpoint on a branch miss.
// Allocate checkpoint on a branch queue

always_ff @(posedge clk)
if (rst) begin
	state <= CHKPT_IDLE;
	alloc_chkpt <= FALSE;
	ialloc_chkpt <= FALSE;
	setcp <= FALSE;
	cndx <= {$bits(checkpt_ndx_t){1'b0}};
	setcp_grp <= 6'd0;
end
else begin
	ialloc_chkpt <= FALSE;
	alloc_chkpt <= FALSE;
	setcp <= FALSE;
	case (state)
	CHKPT_IDLE:
		begin
			if (restore) begin
				$display("Restoring checkpint %d.", miss_cp);
				cndx <= miss_cp;
			end
			for (n1 = 0; n1 < Qupls4_pkg::ROB_ENTRIES/4; n1 = n1 + 1) begin
				if (pgh[n1].v && pgh[n1].has_branch && !pgh[n1].cndxv) begin
					ialloc_chkpt <= TRUE;
					setcp_grp <= n1;
					state <= CHKPT_ALLOC1;
				end
				else if (pgh[n1].v && !pgh[n1].cndxv) begin
					setcp_grp <= n1;
					state <= CHKPT_SET;
				end
			end
		end
	CHKPT_ALLOC1:
		state <= CHKPT_ALLOC2;
	CHKPT_ALLOC2:
		if (!chkpt_stall) begin
			$display("Setting new checkpoint %d.", avail_chkpt[0]);
			alloc_chkpt <= TRUE;
			cndx <= avail_chkpt[0];
			setcp <= TRUE;
			state <= CHKPT_IDLE;
		end
	CHKPT_SET:
		begin
			$display("Setting checkpoint %d.", cndx);
			setcp <= TRUE;
			state <= CHKPT_IDLE;
		end
	endcase
end

reg [3:0] free_chkpt_is;
reg [3:0] free_chkpt2s;
checkpt_ndx_t fchkpt;
checkpt_ndx_t [3:0] fchkpt_is;
checkpt_ndx_t [3:0] fchkpt2s;
always_comb free_chkpt_is[0] = free_chkpt;
always_comb free_chkpt_is[1] = free_chkpt;
always_comb free_chkpt_is[2] = free_chkpt;
always_comb free_chkpt_is[3] = free_chkpt;
always_comb fchkpt_is[0] = fchkpt;
always_comb fchkpt_is[1] = fchkpt;
always_comb fchkpt_is[2] = fchkpt;
always_comb fchkpt_is[3] = fchkpt;
always_comb free_chkpt2s[0] = free_chkpt2;
always_comb free_chkpt2s[1] = free_chkpt2;
always_comb free_chkpt2s[2] = free_chkpt2;
always_comb free_chkpt2s[3] = free_chkpt2;
always_comb fchkpt2s[0] = fchkpt2;
always_comb fchkpt2s[1] = fchkpt2;
always_comb fchkpt2s[2] = fchkpt2;
always_comb fchkpt2s[3] = fchkpt2;

// Checkpoint allocator / deallocator
// GROUP_ALLOC if (TRUE) allocates a single checkpoint for the instruction group.

Qupls4_checkpoint_allocator
#(.GROUP_ALLOC(TRUE))
uchkpta1
(
	.rst(rst),
	.clk(clk),
	.clk5x(clk5x),
	.ph4(ph4),
	.alloc_chkpt(ialloc_chkpt),
	.br(4'h0),
	.chkptn(avail_chkpt),
	.free_chkpt_i(free_chkpt_is),
	.fchkpt_i(fchkpt_is),
	.free_chkpt2(free_chkpt2s),
	.fchkpt2(fchkpt2s),
	.chkpts_to_free(chkpts_to_free),
	.stall(chkpt_stall)
);

// Free branch checkpoints once the branch is done.
/*
Qupls4_checkpoint_freer uchkptfr1
(
	.rst(rst),
	.clk(clk),
	.pgh(pgh),
	.free(free_chkpt),
	.chkpt(fchkpt),
	.chkpt_gndx(freecp_grp)
);
*/
/*
always_ff @(posedge clk)
if (rst) begin
	gndx <= 6'd0;
	free_chkpt2 <= FALSE;
	backout_st2 <= 2'd0;
	grpcnt <= 6'd0;
end
else begin
	free_chkpt2 <= FALSE;
	case(backout_st2)
	2'd0:
		if (restore) begin
			gndx <= ((fcu_id + 3'd4) % Qupls4_pkg::ROB_ENTRIES) >> 2;
			backout_st2 <= 2'd1;
			grpcnt <= 6'd0;
		end
	2'd1:
		begin
			if (pgh[gndx].cndx != pgh[fcu_id>>2].cndx && pgh[gndx].sn > pgh[fcu_id>>2].sn) begin
				free_chkpt2 <= TRUE;
				fchkpt2 <= pgh[gndx].cndx;
			end 
			gndx <= (gndx + 3'd1) % (Qupls4_pkg::ROB_ENTRIES/4);
		end
	endcase
end
*/

endmodule
