// ============================================================================
//        __
//   \\__/ o\    (C) 2023-2025  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
//
// ============================================================================

import const_pkg::*;
import Qupls4_pkg::*;

module Qupls4_info(ndx, coreno, thread, o);
input [63:0] coreno;
input [2:0] thread;
input [4:0] ndx;
output cpu_types_pkg::value_t o;

always_comb
	case(ndx)
	5'd0:	o = coreno;
	5'd1:	o = {61'd0,thread};
	5'd2:	o = "Finitron";
	5'd3:	o = 64'd0;
	5'd4:	o = "64BitSS ";
	5'd5: o = 64'd0;
	5'd6:	o = "Qupls4  ";
	5'd7:	o = 64'd0;
	5'd8:	o = "M1";
	5'd9:	o = 64'h1234;
	5'd10:	o = 64'h0;
	5'd11:	
		begin
			o[31:0] = 32'd32768;
			o[63:32] = 32'd65536;
		end
	5'd12:	o = 64'd8;
	5'd13:	o = 64'd64;
	default:	o = 64'h0;
	endcase
	
endmodule
