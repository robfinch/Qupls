
 	if (ns_dstregv[0][0]) begin rob[ns_rndx_o[0]].op.pRd  <= ns_dstreg[0][0]; rob[ns_rndx_o[0]].op.pRdv <= TRUE; end
 	if (ns_dstregv[0][1]) begin rob[ns_rndx_o[0]].op.pRd2 <= ns_dstreg[0][1]; rob[ns_rndx_o[0]].op.pRd2v <= TRUE; end
 	if (ns_dstregv[0][2]) begin rob[ns_rndx_o[0]].op.pRco <= ns_dstreg[0][2]; rob[ns_rndx_o[0]].op.pRcov <= TRUE; end

 	if (ns_dstregv[1][0]) begin rob[ns_rndx_o[1]].op.pRd  <= ns_dstreg[1][0]; rob[ns_rndx_o[1]].op.pRdv <= TRUE; end
 	if (ns_dstregv[1][1]) begin rob[ns_rndx_o[1]].op.pRd2 <= ns_dstreg[1][1]; rob[ns_rndx_o[1]].op.pRd2v <= TRUE; end
 	if (ns_dstregv[1][2]) begin rob[ns_rndx_o[1]].op.pRco <= ns_dstreg[1][2]; rob[ns_rndx_o[1]].op.pRcov <= TRUE; end

 	if (ns_dstregv[2][0]) begin rob[ns_rndx_o[2]].op.pRd  <= ns_dstreg[2][0]; rob[ns_rndx_o[2]].op.pRdv <= TRUE; end
 	if (ns_dstregv[2][1]) begin rob[ns_rndx_o[2]].op.pRd2 <= ns_dstreg[2][1]; rob[ns_rndx_o[2]].op.pRd2v <= TRUE; end
 	if (ns_dstregv[2][2]) begin rob[ns_rndx_o[2]].op.pRco <= ns_dstreg[2][2]; rob[ns_rndx_o[2]].op.pRcov <= TRUE; end

 	if (ns_dstregv[3][0]) begin rob[ns_rndx_o[3]].op.pRd  <= ns_dstreg[3][0]; rob[ns_rndx_o[3]].op.pRdv <= TRUE; end
 	if (ns_dstregv[3][1]) begin rob[ns_rndx_o[3]].op.pRd2 <= ns_dstreg[3][1]; rob[ns_rndx_o[3]].op.pRd2v <= TRUE; end
 	if (ns_dstregv[3][2]) begin rob[ns_rndx_o[3]].op.pRco <= ns_dstreg[3][2]; rob[ns_rndx_o[3]].op.pRcov <= TRUE; end

