// ============================================================================
//        __
//   \\__/ o\    (C) 2021-2023  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Given a "flat" or unnormalized address, convert it into block,group,and num
// ============================================================================

import QuplsPkg::*;

module Qupls_norm_addr(misspc, ibh, len0, len1, len2, missblock, missgrp, missinsn);
input pc_address_t misspc;	// unnormalized miss address
input ibh_t ibh;						// instruction block header
input [2:0] len0;
input [2:0] len1;
input [2:0] len2;
output reg [$bits(pc_address_t)-1:6] missblock;
output reg [2:0] missgrp;		// group instruction is contained in
output reg [2:0] missinsn;	// instruction number of address

reg [5:0] grpndx;						// byte index of instruction in group

assign missblock = misspc[$bits(pc_address_t)-1:6];

function [2:0] fnInsnNum;
input [5:0] pc;
input [5:0] offs;
reg [5:0] grpndx;
begin
	grpndx = pc - offs;
	// Sort
	if (grpndx > len0+len1+len2)
		fnInsnNum = 3'd3;
	else if (grpndx > len0+len1)
		fnInsnNum = 3'd2;
	else if (grpndx > len0)
		fnInsnNum = 3'd1;
	else
		fnInsnNum = 3'd0;					// assume first instruction
end			
endfunction

always_comb
begin
	if (misspc[5:0] >= ibh.offs[3])
		missgrp = 3'd4;
	else if (misspc[5:0] >= ibh.offs[2])
		missgrp = 3'd3;
	else if (misspc[5:0] >= ibh.offs[1])
		missgrp = 3'd2;
	else if (misspc[5:0] >= ibh.offs[0])
		missgrp = 3'd1;
	else
		missgrp = 3'd0;

	if (missgrp==3'd0)
		missinsn = fnInsnNum(misspc[5:0], ibh.offs[0]);
	else if (missgpr==3'd1)
		missinsn = fnInsnNum(misspc[5:0], ibh.offs[1]);
	else if (missgpr==3'd2)
		missinsn = fnInsnNum(misspc[5:0], ibh.offs[2]);
	else if (missgpr==3'd3)
		missinsn = fnInsnNum(misspc[5:0], ibh.offs[3]);
	else
		missinsn = fnInsnNum(misspc[5:0], ibh.offs[4]);
end

endmodule
