// ============================================================================
//        __
//   \\__/ o\    (C) 2023-2025  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================

import Stark_pkg::*;

module Stark_decode_multicycle(instr, multicycle);
input Stark_pkg::instruction_t instr;
output multicycle;

function fnIsMC;
input Stark_pkg::instruction_t ir;
begin
	case(ir.any.opcode)
	Stark_pkg::OP_FLT:
		case(ir.fpu.op4)
		Stark_pkg::FOP4_FMUL,Stark_pkg::FOP4_FDIV,Stark_pkg::FOP4_FADD,Stark_pkg::FOP4_FSUB:
			fnIsMC = 1'b1;
		Stark_pkg::FOP4_G8:
			case (ir.fpu.op3)
			Stark_pkg::FG8_SCALEB:	fnIsMC = 1'b1;
			default:
				fnIsMC = 1'b0;
			endcase
		Stark_pkg::FOP4_G10:	fnIsMC = 1'b1;
		Stark_pkg::FOP4_TRIG: fnIsMC = 1'b1;
		default:	fnIsMC = 1'b0;
		endcase
	Stark_pkg::OP_MUL:
		fnIsMC = 1'b1;
	Stark_pkg::OP_DIV:
	 	fnIsMC = 1'b1;
	default:	fnIsMC = 1'b0;
	endcase
end
endfunction

assign multicycle = fnIsMC(instr);

endmodule
