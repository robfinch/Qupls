// ============================================================================
//        __
//   \\__/ o\    (C) 2021-2025  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================

import Qupls4_pkg::*;

module Qupls4_decode_sau(instr, sau);
input Qupls4_pkg::micro_op_t instr;
output sau;

function fnIsSau;
input Qupls4_pkg::micro_op_t ir;
begin
	fnIsSau = 1'b0;
	case(ir.opcode)
	Qupls4_pkg::OP_BFLD:
		fnIsSau = 1'b1;
	Qupls4_pkg::OP_R3B,Qupls4_pkg::OP_R3W,Qupls4_pkg::OP_R3T,Qupls4_pkg::OP_R3O,
	Qupls4_pkg::OP_R3BP,Qupls4_pkg::OP_R3WP,Qupls4_pkg::OP_R3TP,Qupls4_pkg::OP_R3OP,
	Qupls4_pkg::OP_R3P:
		fnIsSau = 1'b1;
	Qupls4_pkg::OP_FLTH,Qupls4_pkg::OP_FLTS,Qupls4_pkg::OP_FLTD,Qupls4_pkg::OP_FLTQ,
	Qupls4_pkg::OP_FLTPH,Qupls4_pkg::OP_FLTPS,Qupls4_pkg::OP_FLTPD,Qupls4_pkg::OP_FLTPQ,
	Qupls4_pkg::OP_FLTP:
		case(ir.func)
		Qupls4_pkg::FLT_CMP,
		Qupls4_pkg::FLT_ABS,Qupls4_pkg::FLT_NEG:
			fnIsSau = 1'b1;
		default:	fnIsSau = 1'b0;
		endcase
	Qupls4_pkg::OP_CHK:	fnIsSau = 1'b1;
	Qupls4_pkg::OP_ADDI:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_SUBFI:	fnIsSau = 1'b1;
	Qupls4_pkg::OP_CMPI:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_CMPUI:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_ANDI:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_ORI:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_XORI:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_SHIFT:	fnIsSau = 1'b1;
	Qupls4_pkg::OP_CSR:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_MOVMR:		fnIsSau = 1'b1;
	Qupls4_pkg::OP_LOADA:	fnIsSau = 1'b1;
	Qupls4_pkg::OP_NOP,
	Qupls4_pkg::OP_PUSH,Qupls4_pkg::OP_POP:
		fnIsSau = 1'b1;
	Qupls4_pkg::OP_FENCE:
		fnIsSau = 1'b1;
	default:
		fnIsSau = 1'b0;
	endcase
end
endfunction

assign sau = fnIsSau(instr);

endmodule
