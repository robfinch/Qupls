// ============================================================================
//        __
//   \\__/ o\    (C) 2021-2024  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================

import cpu_types_pkg::*;
import QuplsPkg::*;

module Qupls_decode_Rb(om, ipl, instr, has_immb, Rb, Rbz, Rbn);
input operating_mode_t om;
input [2:0] ipl;
input ex_instruction_t instr;
input has_immb;
output cpu_types_pkg::aregno_t Rb;
output reg Rbz;
output reg Rbn;

function aregno_t fnRb;
input ex_instruction_t ir;
input has_immb;
begin
	case(ir.ins.any.opcode)
	OP_RTD:
		fnRb = 9'd31;
	OP_FLT3:
		fnRb = ir.aRb;
	default:
		if (has_immb)
			fnRb = 9'd0;
		else if (ir.ins.any.opcode==OP_LDX && ir.ins.lsn.func==FN_LDCTX)
			fnRb = 9'd0;
		else if (ir.ins.any.opcode==OP_STX && ir.ins.lsn.func==FN_STCTX)
			fnRb = 9'd0;
		else if (fnImmb(ir))
			fnRb = 9'd0;
		else
			fnRb = ir.aRb;
	endcase
end
endfunction

always_comb
begin
	Rb = fnRb(instr, has_immb);
	if (Rb==9'd31)
		Rb = 9'd32|om;
	Rbn = instr.ins.r3.Rb.n;
	Rbz = ~|Rb;
end

endmodule

